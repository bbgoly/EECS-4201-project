// ----  Probes  ----
`define PROBE_ADDR addr
`define PROBE_DATA_IN data_in
`define PROBE_DATA_OUT data_out
`define PROBE_READ_EN read_en
`define PROBE_WRITE_EN write_en

`define PROBE_F_PC f_pc
`define PROBE_F_INSN f_insn
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd1
// ----  Top module  ----
