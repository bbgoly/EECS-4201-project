// ----  Probes  ----
`define PROBE_F_PC f_pc
`define PROBE_F_INSN f_insn

`define PROBE_D_PC d_pc
`define PROBE_D_OPCODE d_opcode
`define PROBE_D_RD d_rd
`define PROBE_D_FUNCT3 d_funct3
`define PROBE_D_RS1 d_rs1
`define PROBE_D_RS2 d_rs2
`define PROBE_D_FUNCT7 d_funct7
`define PROBE_D_IMM d_imm
`define PROBE_D_SHAMT d_shamt

`define PROBE_R_WRITE_ENABLE r_write_enable
`define PROBE_R_WRITE_DESTINATION r_write_destination
`define PROBE_R_WRITE_DATA r_write_data
`define PROBE_R_READ_RS1 r_read_rs1
`define PROBE_R_READ_RS2 r_read_rs2
`define PROBE_R_READ_RS1_DATA r_read_rs1_data
`define PROBE_R_READ_RS2_DATA r_read_rs2_data

`define PROBE_E_PC e_pc
`define PROBE_E_ALU_RES e_alu_res
`define PROBE_E_BR_TAKEN e_br_taken

// `define PROBE_M_PC                // ??
// `define PROBE_M_ADDRESS           // ??
// `define PROBE_M_SIZE_ENCODED      // ??
// `define PROBE_M_DATA              // ??

// `define PROBE_W_PC                // ??
// `define PROBE_W_ENABLE            // ??
// `define PROBE_W_DESTINATION       // ??
// `define PROBE_W_DATA              // ??
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd4 
// ----  Top module  ----
