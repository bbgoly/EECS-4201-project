/*
 * Yousif Kndkji
 * Salman Kayani
 * Module: writeback
 *
 * Description: Write-back control stage implementation
 *
 * Inputs:
 * 1) PC pc_i
 * 2) result from alu alu_res_i
 * 3) data from memory memory_data_i
 * 4) data to select for write-back wbsel_i
 *
 * Outputs:
 * 1) DWIDTH wide write back data write_data_o
 */

`include "constants.svh"

module writeback #(
    parameter int DWIDTH=32,
    parameter int AWIDTH=32
)(
	input logic [AWIDTH-1:0] pc_i,
	input logic [DWIDTH-1:0] alu_res_i,
	input logic [DWIDTH-1:0] memory_data_i,
	input logic [1:0] wbsel_i,
	// input logic brtaken_i,
	
	output logic [DWIDTH-1:0] writeback_data_o
);

    always_comb begin
        unique case (wbsel_i)
            WB_ALU: writeback_data_o = alu_res_i;      	// R-type, I-type ALU operations
            WB_MEM: writeback_data_o = memory_data_i;  	// Load instructions
            WB_PC: writeback_data_o = pc_i + 32'd4;		// JAL / JALR link return value
            default: writeback_data_o = alu_res_i;		// ALU result as default
        endcase
    end

endmodule : writeback